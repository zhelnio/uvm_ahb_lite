/********************************************************************                                                                                                  
 * Copyright (c) 2014
 * All rights reserved.
 *   
 * \file    ahb_sequence_lib.svh
 * \brief   
 * \version 1.0
 * \author  seabeam
 * \Email   seabeam@sina.com
 * \date    2014-11-29
 ********************************************************************/
`ifndef AHB_CASE_PKG_SV
`define AHB_CASE_PKG_SV
               
package ahb_case_pkg;
    import uvm_pkg::*;
    import ahb_pkg::*;                                                                                                                                                 
                  
    `include "uvm_macros.svh"
               
    `include "ahb_case_base.svh"
endpackage     
               
`endif 
