/********************************************************************
 * Copyright (c) 2014
 * All rights reserved.
 *
 * \file    amba_define.svh
 * \brief   
 * \version 1.0
 * \author  seabeam
 * \Email   seabeam@sina.com
 * \date    2014-12-18
 ********************************************************************/

`ifndef AMBA_DEFINE_SVH
`define AMBA_DEFINE_SVH

    `ifndef AMBA_BUS_DATA_WIDTH
        `define AMBA_BUS_DATA_WIDTH     32
    `endif
    `ifndef AMBA_BUS_ADDR_WIDTH
        `define AMBA_BUS_ADDR_WIDTH     32
    `endif

`endif
